-- SCOMP Interface: Handle Commands + Pulse Logic
PROCESS (RESETN, CS)
    VARIABLE command : STD_LOGIC_VECTOR(3 DOWNTO 0);
    VARIABLE led_index : INTEGER RANGE 0 TO 9;
BEGIN
    IF RESETN = '0' THEN
        led_state <= (OTHERS => '0');
        led_brightness <= (OTHERS => "1111");
        led_gamma <= (OTHERS => '1');
        -- pulse mode variables
        led_pulse_mode <= (OTHERS => '0');
        led_pulse_brightness <= (OTHERS => "0000");
        pulse_clock <= 0;
        led_pulse_flag <= (OTHERS => '0');
        led_pulse_enabled <= (OTHERS => '0');
        led_pulse_target <= (OTHERS => "0000");
        led_pulse_counter <= (OTHERS => 0);

    ELSIF rising_edge(CS) THEN

        -- Handle WRITE commands
        IF WRITE_EN = '1' THEN
            command := IO_DATA(15 DOWNTO 12);
            led_index := CONV_INTEGER(IO_DATA(11 DOWNTO 8));

            CASE command IS
                WHEN "0000" =>  -- F1 Set all LEDs directly
                    led_state <= IO_DATA(9 DOWNTO 0);

                WHEN "0001" =>  -- F2.1 Set individual LED ON
                    IF led_index <= 9 THEN
                        led_state(led_index) <= '1';
                    END IF;

                WHEN "0010" =>  -- F2.2 Clear individual LED
                    IF led_index <= 9 THEN
                        led_state(led_index) <= '0';
                    END IF;

                WHEN "0011" =>  -- F2.3 Toggle individual LED
                    IF led_index <= 9 THEN
                        led_state(led_index) <= NOT led_state(led_index);
                    END IF;

                WHEN "0100" =>  -- F3 Set individual brightness + gamma
                    IF led_index <= 9 THEN
                        led_brightness(led_index) <= IO_DATA(3 DOWNTO 0);
                        led_gamma(led_index) <= IO_DATA(4);
                        led_state(led_index) <= '1';
                    END IF;

                WHEN "0101" =>  -- F4 Set all brightness + gamma
                    FOR i IN 0 TO 9 LOOP
                        led_brightness(i) <= IO_DATA(3 DOWNTO 0);
                        led_gamma(i) <= IO_DATA(4);
                        led_state(i) <= '1';
                    END LOOP;

                WHEN "0111" =>  -- F7: Individual pulse mode
                    IF led_index <= 9 THEN
                        led_pulse_enabled(led_index) <= '1';
                        led_pulse_target(led_index) <= IO_DATA(3 DOWNTO 0);
                        led_pulse_counter(led_index) <= 0;
                    END IF;

                WHEN "1010" =>  -- F8: ripple mode
                    ripple_mode <= '1';

                WHEN OTHERS =>
                    NULL;
            END CASE;
        END IF;

        -- Commented legacy pulse logic
        -- IF pulse_mode = '1' AND command = "0111" THEN
        --     IF pulse_clock < 74999 THEN
        --         pulse_clock <= pulse_clock + 1;
        --     ELSE
        --         pulse_clock <= 0;
        --         IF pulse_flag = '0' THEN
        --             -- We're in the increasing phase
        --             IF pulse_brightness = "1111" THEN
        --                 pulse_flag <= '1';
        --                 pulse_brightness <= pulse_brightness - 1;
        --             ELSE
        --                 pulse_brightness <= pulse_brightness + 1;
        --             END IF;
        --         ELSE
        --             -- We're in the decreasing phase
        --             IF pulse_brightness = "0000" THEN
        --                 pulse_flag <= '0';
        --                 pulse_brightness <= pulse_brightness + 1;
        --             ELSE
        --                 pulse_brightness <= pulse_brightness - 1;
        --             END IF;
        --         END IF;
        --     END IF;
        -- END IF;

        -- Update all LEDs with current brightness
        FOR i IN 0 TO 9 LOOP
            IF led_pulse_enabled(i) = '1' THEN
                IF led_pulse_counter(i) < (37500 * (CONV_INTEGER(led_pulse_target(i)) + 1)) THEN
                    led_pulse_counter(i) <= led_pulse_counter(i) + 1;
                ELSE
                    led_pulse_counter(i) <= 0;
                    IF led_pulse_flag(i) = '0' THEN
                        -- We're in the increasing phase
                        IF led_pulse_brightness(i) = "1111" THEN
                            led_pulse_flag(i) <= '1';
                            led_pulse_brightness(i) <= led_pulse_brightness(i) - 1;
                        ELSE
                            led_pulse_brightness(i) <= led_pulse_brightness(i) + 1;
                        END IF;
                    ELSE
                        -- We're in the decreasing phase
                        IF led_pulse_brightness(i) = "0000" THEN
                            led_pulse_flag(i) <= '0';
                            led_pulse_brightness(i) <= led_pulse_brightness(i) + 1;
                        ELSE
                            led_pulse_brightness(i) <= led_pulse_brightness(i) - 1;
                        END IF;
                    END IF;
                    led_gamma(i) <= '1';
                    led_state(i) <= '1';
                END IF;
            END IF;
        END LOOP;

    END IF;
END PROCESS;